--=============================
-- Listing 9.1 async clear
--=============================
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity mod10_counter is
   port(
      clk, reset: in std_logic;
      q: out std_logic_vector(3 downto 0)
   );
end mod10_counter;
 
--architecture poor_async_arch of mod10_counter is
--   signal r_reg: unsigned(3 downto 0);
--   signal r_next: unsigned(3 downto 0);
--   signal async_clr: std_logic;
--begin
--   -- register
--   process(clk,async_clr)
--   begin
--      if (async_clr='1') then
--         r_reg <= (others=>'0');
--      elsif (clk'event and clk='1') then
--         r_reg <= r_next;
--      end if;
--   end process;
--   -- asynchronous clear
--   async_clr <= '1' when (reset='1' or r_reg="1010") else
--                '0';
--   -- next state logic
--   r_next <= r_reg + 1;
--   -- output logic
--   q <= std_logic_vector(r_reg);
--end poor_async_arch;
-- 
 
--=============================
-- Listing 9.2
--=============================
architecture two_seg_arch of mod10_counter is
   signal r_reg: unsigned(3 downto 0);
   signal r_next: unsigned(3 downto 0);
begin
   -- register
   process(clk,reset)
   begin
      if (reset='1') then
         r_reg <= (others=>'0');
      elsif (clk'event and clk='1') then
         r_reg <= r_next;
      end if;
   end process;
   -- next-state logic
   r_next <= (others=>'0') when r_reg=9 else
             r_reg + 1;
   -- output logic
   q <= std_logic_vector(r_reg);
end two_seg_arch;