--=============================
-- Listing 9.3 gated clock
--=============================
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity binary_counter is
   port(
      clk, reset: in std_logic;
      en: in std_logic;
      q: out std_logic_vector(3 downto 0)
   );
end binary_counter;

--architecture gated_clk_arch of binary_counter is
--   signal r_reg: unsigned(3 downto 0);
--   signal r_next: unsigned(3 downto 0);
--   signal gated_clk: std_logic;
--begin
--   -- register
--   process(gated_clk,reset)
--   begin
--      if (reset='1') then
--         r_reg <= (others=>'0');
--      elsif (gated_clk'event and gated_clk='1') then
--         r_reg <= r_next;
--      end if;
--   end process;
--   -- gated clock
--   gated_clk <= clk and en;
--   -- next-state logic
--   r_next <= r_reg + 1;
--   -- output logic
--   q <= std_logic_vector(r_reg);
--end gated_clk_arch;

--=============================
-- Listing 9.4
--=============================
architecture two_seg_arch of binary_counter is
   signal r_reg: unsigned(3 downto 0);
   signal r_next: unsigned(3 downto 0);
begin
   -- register
   process(clk,reset)
   begin
      if (reset='1') then
         r_reg <= (others=>'0');
      elsif (clk'event and clk='1') then
         r_reg <= r_next;
      end if;
   end process;
   -- next-state logic
   r_next <= r_reg + 1 when en='1' else
             r_reg;
   -- output logic
   q <= std_logic_vector(r_reg);
end two_seg_arch;